module simple_display();

  initial begin
    $display("\n\t Write your Message here");
  end

endmodule